package bus_pkg;
  `include "dBus_if.sv"
  `include "iBus_if.sv"
  `include "intrBus_if.sv"
  `include "debug_if.sv"
endpackage
