typedef uvm_sequencer#(ibus_tx) ibus_sqr;
