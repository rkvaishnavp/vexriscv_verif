class dbus_tx extends uvm_sequence_item;

  int 

  function new(string name = "dbus_tx");
    super.new(name);
  endfunction //new()
endclass //dbus_tx extends uvm_sequence_item