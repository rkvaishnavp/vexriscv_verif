typedef uvm_sequencer#(dbus_tx) dbus_sqr;
