class VexRiscv_cov extends uvm_coverage;
  function new();
    
  endfunction //new()
endclass //VexRiscv_cov extends uvm_coverage