typedef uvm_sequencer#(debug_tx) debug_sqr;
